module Statistics_8Bin(
  input                   iclk,
  input                   ireset,
  input         [17:0]    igradient0,
  input         [17:0]    igradient1,
  input         [17:0]    igradient2,
  input         [17:0]    igradient3,
  input         [17:0]    igradient4,
  input         [17:0]    igradient5,
  input         [17:0]    igradient6,
  input         [17:0]    igradient7,
  input         [17:0]    igradient8,
  input         [17:0]    igradient9,
  input         [17:0]    igradient10,
  input         [17:0]    igradient11,
  input         [17:0]    igradient12,
  input         [17:0]    igradient13,
  input         [17:0]    igradient14,
  input         [17:0]    igradient15,
  output        [12:0]    obin_value0,
  output        [12:0]    obin_value1,
  output        [12:0]    obin_value2,
  output        [12:0]    obin_value3,
  output        [12:0]    obin_value4,
  output        [12:0]    obin_value5,
  output        [12:0]    obin_value6,
  output        [12:0]    obin_value7
);

StatisticsBin Statistics_8Bin1(
  .iclk(iclk),
  .ireset(ireset),
  .iline0(igradient0),
  .iline1(igradient1),
  .iline2(igradient2),
  .iline3(igradient3),
  .iline4(igradient4),
  .iline5(igradient5),
  .iline6(igradient6),
  .iline7(igradient7),
  .iline8(igradient8),
  .iline9(igradient9),
  .iline10(igradient10),
  .iline11(igradient11),
  .iline12(igradient12),
  .iline13(igradient13),
  .iline14(igradient14),
  .iline15(igradient15),
  .ilower_limit(9'd0),
  .iupper_limit(9'd45),
  .obin_value(obin_value0)
);

StatisticsBin Statistics_8Bin2(
  .iclk(iclk),
  .ireset(ireset),
  .iline0(igradient0),
  .iline1(igradient1),
  .iline2(igradient2),
  .iline3(igradient3),
  .iline4(igradient4),
  .iline5(igradient5),
  .iline6(igradient6),
  .iline7(igradient7),
  .iline8(igradient8),
  .iline9(igradient9),
  .iline10(igradient10),
  .iline11(igradient11),
  .iline12(igradient12),
  .iline13(igradient13),
  .iline14(igradient14),
  .iline15(igradient15),
  .ilower_limit(9'd45),
  .iupper_limit(9'd90),
  .obin_value(obin_value1)
);

StatisticsBin Statistics_8Bin3(
  .iclk(iclk),
  .ireset(ireset),
  .iline0(igradient0),
  .iline1(igradient1),
  .iline2(igradient2),
  .iline3(igradient3),
  .iline4(igradient4),
  .iline5(igradient5),
  .iline6(igradient6),
  .iline7(igradient7),
  .iline8(igradient8),
  .iline9(igradient9),
  .iline10(igradient10),
  .iline11(igradient11),
  .iline12(igradient12),
  .iline13(igradient13),
  .iline14(igradient14),
  .iline15(igradient15),
  .ilower_limit(9'd90),
  .iupper_limit(9'd135),
  .obin_value(obin_value2)
);

StatisticsBin Statistics_8Bin4(
  .iclk(iclk),
  .ireset(ireset),
  .iline0(igradient0),
  .iline1(igradient1),
  .iline2(igradient2),
  .iline3(igradient3),
  .iline4(igradient4),
  .iline5(igradient5),
  .iline6(igradient6),
  .iline7(igradient7),
  .iline8(igradient8),
  .iline9(igradient9),
  .iline10(igradient10),
  .iline11(igradient11),
  .iline12(igradient12),
  .iline13(igradient13),
  .iline14(igradient14),
  .iline15(igradient15),
  .ilower_limit(9'd135),
  .iupper_limit(9'd180),
  .obin_value(obin_value3)
);

StatisticsBin Statistics_8Bin5(
  .iclk(iclk),
  .ireset(ireset),
  .iline0(igradient0),
  .iline1(igradient1),
  .iline2(igradient2),
  .iline3(igradient3),
  .iline4(igradient4),
  .iline5(igradient5),
  .iline6(igradient6),
  .iline7(igradient7),
  .iline8(igradient8),
  .iline9(igradient9),
  .iline10(igradient10),
  .iline11(igradient11),
  .iline12(igradient12),
  .iline13(igradient13),
  .iline14(igradient14),
  .iline15(igradient15),
  .ilower_limit(9'd180),
  .iupper_limit(9'd225),
  .obin_value(obin_value4)
);

StatisticsBin Statistics_8Bin6(
  .iclk(iclk),
  .ireset(ireset),
  .iline0(igradient0),
  .iline1(igradient1),
  .iline2(igradient2),
  .iline3(igradient3),
  .iline4(igradient4),
  .iline5(igradient5),
  .iline6(igradient6),
  .iline7(igradient7),
  .iline8(igradient8),
  .iline9(igradient9),
  .iline10(igradient10),
  .iline11(igradient11),
  .iline12(igradient12),
  .iline13(igradient13),
  .iline14(igradient14),
  .iline15(igradient15),
  .ilower_limit(9'd225),
  .iupper_limit(9'd270),
  .obin_value(obin_value5)
);

StatisticsBin Statistics_8Bin7(
  .iclk(iclk),
  .ireset(ireset),
  .iline0(igradient0),
  .iline1(igradient1),
  .iline2(igradient2),
  .iline3(igradient3),
  .iline4(igradient4),
  .iline5(igradient5),
  .iline6(igradient6),
  .iline7(igradient7),
  .iline8(igradient8),
  .iline9(igradient9),
  .iline10(igradient10),
  .iline11(igradient11),
  .iline12(igradient12),
  .iline13(igradient13),
  .iline14(igradient14),
  .iline15(igradient15),
  .ilower_limit(9'd270),
  .iupper_limit(9'd315),
  .obin_value(obin_value6)
);

StatisticsBin Statistics_8Bin8(
  .iclk(iclk),
  .ireset(ireset),
  .iline0(igradient0),
  .iline1(igradient1),
  .iline2(igradient2),
  .iline3(igradient3),
  .iline4(igradient4),
  .iline5(igradient5),
  .iline6(igradient6),
  .iline7(igradient7),
  .iline8(igradient8),
  .iline9(igradient9),
  .iline10(igradient10),
  .iline11(igradient11),
  .iline12(igradient12),
  .iline13(igradient13),
  .iline14(igradient14),
  .iline15(igradient15),
  .ilower_limit(9'd315),
  .iupper_limit(9'd360),
  .obin_value(obin_value7)
);

endmodule 